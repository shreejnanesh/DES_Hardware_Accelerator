
package enc_pkg;

	import uvm_pkg::*;
	`include "grDesEnc.sv"
	`include "sequenceItem.sv"
	`include "driver.sv"
	`include "sequence.sv"
	`include "monitor.sv"
	`include "scoreboard.sv"
	`include "subscriber.sv"
	`include "agent.sv"
	`include "environment.sv"
	`include "test.sv"

endpackage